`define Q0_LN0
`define Q0_LN0_PMA_WIDTH 20
`define Q0_LN0_TX_GEARBOX 1
`define Q0_LN0_RX_GEARBOX 1
`define Q0_LN0_CHANNEL_BONDING_MASTER_SEL 0
`define Q0_LN0_TX_IF_MST_SEL 0
`define Q0_LN1
`define Q0_LN1_PMA_WIDTH 20
`define Q0_LN1_TX_GEARBOX 1
`define Q0_LN1_RX_GEARBOX 1
`define Q0_LN1_CHANNEL_BONDING_MASTER_SEL 0
`define Q0_LN1_TX_IF_MST_SEL 0
`define Q0_LN2
`define Q0_LN2_PMA_WIDTH 20
`define Q0_LN2_TX_GEARBOX 1
`define Q0_LN2_RX_GEARBOX 1
`define Q0_LN2_CHANNEL_BONDING_MASTER_SEL 0
`define Q0_LN2_TX_IF_MST_SEL 0
`define Q0_LN3
`define Q0_LN3_PMA_WIDTH 20
`define Q0_LN3_TX_GEARBOX 1
`define Q0_LN3_RX_GEARBOX 1
`define Q0_LN3_CHANNEL_BONDING_MASTER_SEL 0
`define Q0_LN3_TX_IF_MST_SEL 0
`define MODULE_NAME Customized_PHY_Top
