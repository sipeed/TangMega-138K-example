parameter DRP_NUM = 8;
