`define module_name uart_core
