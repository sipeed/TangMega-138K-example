module color_bar(
	input                 clk,           //pixel clock
	input                 rst,           //reset signal high active

	// output reg [9:0] active_x,              //video x position 
	// output reg [9:0] active_y,             //video y position 

	output                hs,            //horizontal synchronization
	output                vs,            //vertical synchronization
	output                de

);
//     reg         [15:0]  PixelCount;
//     reg         [15:0]  LineCount;

// 	localparam      V_BackPorch = 16'd0; //6
// 	localparam      V_Pluse 	= 16'd5; 
// 	localparam      HightPixel  = 16'd480;
// 	localparam      V_FrontPorch= 16'd45; //62

// 	localparam      H_BackPorch = 16'd182; 	//NOTE: 高像素时钟时，增加这里的延迟，方便K210加入中断
// 	localparam      H_Pluse 	= 16'd1; 
// 	localparam      WidthPixel  = 16'd800; 
// 	localparam      H_FrontPorch= 16'd210;
// endmodule

//800x480
parameter H_ACTIVE = 16'd800;
parameter H_FP = 16'd210;       
parameter H_SYNC = 16'd1;    
parameter H_BP = 16'd182;       
parameter V_ACTIVE = 16'd480; 
parameter V_FP  = 16'd45;     
parameter V_SYNC  = 16'd1;   
parameter V_BP  = 16'd8;     
parameter HS_POL = 1'b0;
parameter VS_POL = 1'b0;

parameter H_TOTAL = H_ACTIVE + H_FP + H_SYNC + H_BP;//horizontal total time (pixels)
parameter V_TOTAL = V_ACTIVE + V_FP + V_SYNC + V_BP;//vertical total time (lines)

reg hs_reg;                      //horizontal sync register
reg vs_reg;                      //vertical sync register
reg[15:0] h_cnt;                 //horizontal counter
reg[15:0] v_cnt;                 //vertical counter
reg h_active;                    //horizontal video active
reg v_active;                    //vertical video active
wire video_active;               //video active(horizontal active and vertical active)
assign hs = hs_reg;
assign vs = vs_reg;

assign de =  h_active & v_active;

always@(posedge clk or posedge rst)
begin
	if(rst == 1'b1)
		h_cnt <= 16'd0;
	else if(h_cnt == H_TOTAL - 1)//horizontal counter maximum value
		h_cnt <= 16'd0;
	else
		h_cnt <= h_cnt + 16'd1;
end

always@(posedge clk or posedge rst)
begin
	if(rst == 1'b1)
		v_cnt <= 16'd0;
	else if(h_cnt == H_FP  - 1)//horizontal sync time
		if(v_cnt == V_TOTAL - 1)//vertical counter maximum value
			v_cnt <= 16'd0;
		else
			v_cnt <= v_cnt + 16'd1;
	else
		v_cnt <= v_cnt;
end

always@(posedge clk or posedge rst)
begin
	if(rst == 1'b1)
		hs_reg <= 1'b0;
	else if(h_cnt == H_FP - 1)//horizontal sync begin
		hs_reg <= HS_POL;
	else if(h_cnt == H_FP + H_SYNC - 1)//horizontal sync end
		hs_reg <= ~hs_reg;
	else
		hs_reg <= hs_reg;
end

always@(posedge clk or posedge rst)
begin
	if(rst == 1'b1)
		h_active <= 1'b0;
	else if(h_cnt == H_FP + H_SYNC + H_BP - 1)//horizontal active begin
		h_active <= 1'b1;
	else if(h_cnt == H_TOTAL - 1)//horizontal active end
		h_active <= 1'b0;
	else
		h_active <= h_active;
end

always@(posedge clk or posedge rst)
begin
	if(rst == 1'b1)
		vs_reg <= 1'd0;
	else if((v_cnt == V_ACTIVE + V_FP + V_SYNC + V_BP) && (h_cnt == H_FP - 1))//vertical sync begin
		vs_reg <= VS_POL;
	else if((v_cnt == V_SYNC) && (h_cnt == H_FP - 1))//vertical sync end
		vs_reg <= ~VS_POL;  
	else
		vs_reg <= vs_reg;
end

always@(posedge clk or posedge rst)
begin
	if(rst == 1'b1)
		v_active <= 1'd0;
	else if((v_cnt == V_SYNC + V_BP) && (h_cnt == H_FP - 1))//vertical active begin
		v_active <= 1'b1;
	else if((v_cnt == V_SYNC + V_BP + V_ACTIVE) && (h_cnt == H_FP - 1)) //vertical active end
		v_active <= 1'b0;   
	else
		v_active <= v_active;
end

endmodule 
